
module ram(clk,rst,in,out);
           input clk;
           input rst;
           input[31:0]in;
           output[31:0]out;
           assign out= in;
           reg xx;
endmodule




